library verilog;
use verilog.vl_types.all;
entity Compare_add_circuit_vlg_vec_tst is
end Compare_add_circuit_vlg_vec_tst;
