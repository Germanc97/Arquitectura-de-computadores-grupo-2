library verilog;
use verilog.vl_types.all;
entity multiplex_vlg_vec_tst is
end multiplex_vlg_vec_tst;
