library verilog;
use verilog.vl_types.all;
entity lab_v1_vlg_check_tst is
    port(
        a               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab_v1_vlg_check_tst;
