library verilog;
use verilog.vl_types.all;
entity lab_v1 is
    port(
        l               : in     vl_logic;
        s               : in     vl_logic;
        d               : in     vl_logic;
        a               : out    vl_logic
    );
end lab_v1;
