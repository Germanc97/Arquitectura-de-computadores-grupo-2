library verilog;
use verilog.vl_types.all;
entity Decoder_vlg_check_tst is
    port(
        salida1         : in     vl_logic;
        salida2         : in     vl_logic;
        salida3         : in     vl_logic;
        salida4         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Decoder_vlg_check_tst;
