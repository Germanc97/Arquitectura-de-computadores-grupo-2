library verilog;
use verilog.vl_types.all;
entity lab_v1_vlg_vec_tst is
end lab_v1_vlg_vec_tst;
