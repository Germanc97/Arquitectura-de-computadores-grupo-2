library verilog;
use verilog.vl_types.all;
entity ram_v1_vlg_vec_tst is
end ram_v1_vlg_vec_tst;
